`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:10:11 01/04/2021 
// Design Name: 
// Module Name:    song 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module song(
	input clk50m,
	input SW,
	output buzzer//high_7s,med_7s,low_7s
    );

//wire [31:0] clkdiv;
//clkdiv divide(clk, clkdiv);
reg speaker;
assign buzzer = SW ? speaker:1'b1;
//output[6:0] high_7s;
//output[6:0] med_7s;
//output[6:0] low_7s;
reg clk_6mhz;
reg clk_4hz;
reg[13:0] divider,origin; reg carry;
reg[10:0] counter; reg[3:0] high,med,low;
reg[2:0] count8;reg[19:0] count20;
always @(posedge clk50m)
    begin if(count8==7) begin count8<=0;clk_6mhz<=1;end
	     else begin count8<=count8+1;clk_6mhz<=0;end
end
always @(posedge clk_6mhz)
    begin
	     if(count20==781250)
		      begin clk_4hz<=~clk_4hz;count20<=0; end
			else  count20<=count20+1;
	end
always @(posedge clk_6mhz)
    begin  if(divider==16383)
	        begin carry<=1;divider<=origin;end
			  else begin divider<=divider+1;carry<=0; end
end
always @(posedge carry)
begin  speaker<=~speaker;end
always @(posedge clk_4hz)
 begin case({high,med,low})
 'h001: origin<=4915;
 'h002: origin<=6168;
 'h003: origin<=7281;
 'h004: origin<=7792;
 'h005: origin<=8730;
 'h006: origin<=9565;
 'h007: origin<=10310;
 'h010: origin<=10647;
 'h020: origin<=11272;
 'h030: origin<=11831;
 'h040: origin<=12094;
 'h050: origin<=12556;
 'h060: origin<=12974;
 'h070: origin<=13346;
 'h100: origin<=13516;
 'h200: origin<=13829;
 'h300: origin<=14109;
 'h400: origin<=14235;
 'h500: origin<=14470;
 'h600: origin<=14678;
 'h700: origin<=14864;
 'h000: origin<=16383;
endcase
end
always @(posedge clk_4hz)
begin
if(counter == 1503) counter<=0;
else counter<=counter+1;
case(counter)
//1
0 :  {high,med,low}<='h020;
1 :  {high,med,low}<='h020;
2 :  {high,med,low}<='h030;
3 :  {high,med,low}<='h030;
4 :  {high,med,low}<='h050;
5 :  {high,med,low}<='h050;
6 :  {high,med,low}<='h010;
7 :  {high,med,low}<='h010;
8 :  {high,med,low}<='h020;
9 :  {high,med,low}<='h020;
10 :  {high,med,low}<='h030;
11 :  {high,med,low}<='h030;
12 :  {high,med,low}<='h050;
13 :  {high,med,low}<='h050;
14 :  {high,med,low}<='h010;
15 :  {high,med,low}<='h010;
//2
16 :  {high,med,low}<='h020;
17 :  {high,med,low}<='h020;
18 :  {high,med,low}<='h030;
19 :  {high,med,low}<='h030;
20 :  {high,med,low}<='h050;
21 :  {high,med,low}<='h050;
22 :  {high,med,low}<='h060;
23 :  {high,med,low}<='h060;
24 :  {high,med,low}<='h020;
25 :  {high,med,low}<='h020;
26 :  {high,med,low}<='h030;
27 :  {high,med,low}<='h030;
28 :  {high,med,low}<='h006;
29 :  {high,med,low}<='h006;
30 :  {high,med,low}<='h010;
31 :  {high,med,low}<='h010;
//3
32 :  {high,med,low}<='h020;
33 :  {high,med,low}<='h020;
34 :  {high,med,low}<='h030;
35 :  {high,med,low}<='h030;
36 :  {high,med,low}<='h050;
37 :  {high,med,low}<='h050;
38 :  {high,med,low}<='h010;
39 :  {high,med,low}<='h010;
40 :  {high,med,low}<='h020;
41 :  {high,med,low}<='h020;
42 :  {high,med,low}<='h030;
43 :  {high,med,low}<='h030;
44 :  {high,med,low}<='h050;
45 :  {high,med,low}<='h050;
46 :  {high,med,low}<='h010;
47 :  {high,med,low}<='h010;
//4
48 :  {high,med,low}<='h020;
49 :  {high,med,low}<='h020;
50 :  {high,med,low}<='h030;
51 :  {high,med,low}<='h030;
52 :  {high,med,low}<='h050;
53 :  {high,med,low}<='h050;
54 :  {high,med,low}<='h060;
55 :  {high,med,low}<='h060;
56 :  {high,med,low}<='h020;
57 :  {high,med,low}<='h020;
58 :  {high,med,low}<='h030;
59 :  {high,med,low}<='h030;
60 :  {high,med,low}<='h006;
61 :  {high,med,low}<='h006;
62 :  {high,med,low}<='h010;
63 :  {high,med,low}<='h010;
//5
64 :  {high,med,low}<='h020;
65 :  {high,med,low}<='h020;
66 :  {high,med,low}<='h030;
67 :  {high,med,low}<='h030;
68 :  {high,med,low}<='h050;
69 :  {high,med,low}<='h050;
70 :  {high,med,low}<='h010;
71 :  {high,med,low}<='h010;
72 :  {high,med,low}<='h020;
73 :  {high,med,low}<='h020;
74 :  {high,med,low}<='h030;
75 :  {high,med,low}<='h030;
76 :  {high,med,low}<='h050;
77 :  {high,med,low}<='h050;
78 :  {high,med,low}<='h010;
79 :  {high,med,low}<='h010;
//6
80 :  {high,med,low}<='h020;
81 :  {high,med,low}<='h020;
82 :  {high,med,low}<='h030;
83 :  {high,med,low}<='h030;
84 :  {high,med,low}<='h050;
85 :  {high,med,low}<='h050;
86 :  {high,med,low}<='h060;
87 :  {high,med,low}<='h060;
88 :  {high,med,low}<='h020;
89 :  {high,med,low}<='h020;
90 :  {high,med,low}<='h030;
91 :  {high,med,low}<='h030;
92 :  {high,med,low}<='h003;
93 :  {high,med,low}<='h003;
94 :  {high,med,low}<='h005;
95 :  {high,med,low}<='h005;
//7
96 :  {high,med,low}<='h006;
97 :  {high,med,low}<='h006;
98 :  {high,med,low}<='h006;
99 :  {high,med,low}<='h006;
100 :  {high,med,low}<='h010;
101 :  {high,med,low}<='h010;
102 :  {high,med,low}<='h020;
103 :  {high,med,low}<='h020;
104 :  {high,med,low}<='h020;
105 :  {high,med,low}<='h020;
106 :  {high,med,low}<='h010;
107 :  {high,med,low}<='h010;
108 :  {high,med,low}<='h005;
109 :  {high,med,low}<='h005;
110 :  {high,med,low}<='h004;
111 :  {high,med,low}<='h004;
//8
112 :  {high,med,low}<='h003;
113 :  {high,med,low}<='h003;
114 :  {high,med,low}<='h005;
115 :  {high,med,low}<='h006;
116 :  {high,med,low}<='h010;
117 :  {high,med,low}<='h010;
118 :  {high,med,low}<='h010;
119 :  {high,med,low}<='h010;
120 :  {high,med,low}<='h000;
121 :  {high,med,low}<='h000;
122 :  {high,med,low}<='h000;
123 :  {high,med,low}<='h000;
124 :  {high,med,low}<='h010;
125 :  {high,med,low}<='h010;
126 :  {high,med,low}<='h007;
127 :  {high,med,low}<='h007;
//9
128 :  {high,med,low}<='h006;
129 :  {high,med,low}<='h006;
130 :  {high,med,low}<='h006;
131 :  {high,med,low}<='h006;
132 :  {high,med,low}<='h010;
133 :  {high,med,low}<='h010;
134 :  {high,med,low}<='h010;
135 :  {high,med,low}<='h010;
136 :  {high,med,low}<='h007;
137 :  {high,med,low}<='h007;
138 :  {high,med,low}<='h005;
139 :  {high,med,low}<='h005;
140 :  {high,med,low}<='h005;
141 :  {high,med,low}<='h005;
142 :  {high,med,low}<='h000;
143 :  {high,med,low}<='h000;
//10
144 :  {high,med,low}<='h005;
145 :  {high,med,low}<='h005;
146 :  {high,med,low}<='h005;
147 :  {high,med,low}<='h005;
148 :  {high,med,low}<='h000;
149 :  {high,med,low}<='h000;
150 :  {high,med,low}<='h000;
151 :  {high,med,low}<='h000;
152 :  {high,med,low}<='h000;
153 :  {high,med,low}<='h000;
154 :  {high,med,low}<='h000;
155 :  {high,med,low}<='h000;
156 :  {high,med,low}<='h003;
157 :  {high,med,low}<='h003;
158 :  {high,med,low}<='h005;
159 :  {high,med,low}<='h005;
//11
160 :  {high,med,low}<='h006;
161 :  {high,med,low}<='h006;
162 :  {high,med,low}<='h006;
163 :  {high,med,low}<='h006;
164 :  {high,med,low}<='h010;
165 :  {high,med,low}<='h010;
166 :  {high,med,low}<='h020;
167 :  {high,med,low}<='h020;
168 :  {high,med,low}<='h020;
169 :  {high,med,low}<='h020;
170 :  {high,med,low}<='h010;
171 :  {high,med,low}<='h010;
172 :  {high,med,low}<='h005;
173 :  {high,med,low}<='h005;
174 :  {high,med,low}<='h004;
175 :  {high,med,low}<='h004;
//12
176 :  {high,med,low}<='h003;
177 :  {high,med,low}<='h003;
178 :  {high,med,low}<='h005;
179 :  {high,med,low}<='h005;
180 :  {high,med,low}<='h007;
181 :  {high,med,low}<='h007;
182 :  {high,med,low}<='h010;
183 :  {high,med,low}<='h010;
184 :  {high,med,low}<='h000;
185 :  {high,med,low}<='h000;
186 :  {high,med,low}<='h000;
187 :  {high,med,low}<='h000;
188 :  {high,med,low}<='h010;
189 :  {high,med,low}<='h010;
190 :  {high,med,low}<='h007;
191 :  {high,med,low}<='h007;
//13
192 :  {high,med,low}<='h006;
193 :  {high,med,low}<='h006;
194 :  {high,med,low}<='h006;
195 :  {high,med,low}<='h006;
196 :  {high,med,low}<='h010;
197 :  {high,med,low}<='h010;
198 :  {high,med,low}<='h010;
199 :  {high,med,low}<='h010;
200 :  {high,med,low}<='h007;
201 :  {high,med,low}<='h007;
202 :  {high,med,low}<='h005;
203 :  {high,med,low}<='h005;
204 :  {high,med,low}<='h000;
205 :  {high,med,low}<='h000;
206 :  {high,med,low}<='h005;
207 :  {high,med,low}<='h005;
//14
208 :  {high,med,low}<='h006;
209 :  {high,med,low}<='h006;
210 :  {high,med,low}<='h006;
211 :  {high,med,low}<='h006;
212 :  {high,med,low}<='h000;
213 :  {high,med,low}<='h000;
214 :  {high,med,low}<='h000;
215 :  {high,med,low}<='h000;
216 :  {high,med,low}<='h000;
217 :  {high,med,low}<='h000;
218 :  {high,med,low}<='h000;
219 :  {high,med,low}<='h000;
220 :  {high,med,low}<='h006;
221 :  {high,med,low}<='h006;
222 :  {high,med,low}<='h007;
223 :  {high,med,low}<='h007;
//15
224 :  {high,med,low}<='h001;
225 :  {high,med,low}<='h001;
226 :  {high,med,low}<='h001;
227 :  {high,med,low}<='h001;
228 :  {high,med,low}<='h001;
229 :  {high,med,low}<='h001;
230 :  {high,med,low}<='h007;
231 :  {high,med,low}<='h007;
232 :  {high,med,low}<='h006;
233 :  {high,med,low}<='h006;
234 :  {high,med,low}<='h007;
235 :  {high,med,low}<='h007;
236 :  {high,med,low}<='h001;
237 :  {high,med,low}<='h001;
238 :  {high,med,low}<='h001;
239 :  {high,med,low}<='h001;
//16
240 :  {high,med,low}<='h000;
241 :  {high,med,low}<='h000;
242 :  {high,med,low}<='h007;
243 :  {high,med,low}<='h007;
244 :  {high,med,low}<='h006;
245 :  {high,med,low}<='h006;
246 :  {high,med,low}<='h007;
247 :  {high,med,low}<='h007;
248 :  {high,med,low}<='h010;
249 :  {high,med,low}<='h010;
250 :  {high,med,low}<='h007;
251 :  {high,med,low}<='h007;
252 :  {high,med,low}<='h005;
253 :  {high,med,low}<='h005;
254 :  {high,med,low}<='h006;
255 :  {high,med,low}<='h006;
//17
256 :  {high,med,low}<='h005;
257 :  {high,med,low}<='h005;
258 :  {high,med,low}<='h001;
259 :  {high,med,low}<='h000;
260 :  {high,med,low}<='h001;
261 :  {high,med,low}<='h001;
262 :  {high,med,low}<='h006;
263 :  {high,med,low}<='h006;
264 :  {high,med,low}<='h005;
265 :  {high,med,low}<='h005;
266 :  {high,med,low}<='h001;
267 :  {high,med,low}<='h001;
268 :  {high,med,low}<='h000;
269 :  {high,med,low}<='h000;
270 :  {high,med,low}<='h002;
271 :  {high,med,low}<='h002;
//18
272 :  {high,med,low}<='h003;
273 :  {high,med,low}<='h003;
274 :  {high,med,low}<='h003;
275 :  {high,med,low}<='h003;
276 :  {high,med,low}<='h000;
277 :  {high,med,low}<='h000;
278 :  {high,med,low}<='h000;
279 :  {high,med,low}<='h000;
280 :  {high,med,low}<='h000;
281 :  {high,med,low}<='h000;
282 :  {high,med,low}<='h000;
283 :  {high,med,low}<='h000;
284 :  {high,med,low}<='h006;
285 :  {high,med,low}<='h006;
286 :  {high,med,low}<='h007;
287 :  {high,med,low}<='h007;
//19
288 :  {high,med,low}<='h010;
289 :  {high,med,low}<='h010;
290 :  {high,med,low}<='h010;
291 :  {high,med,low}<='h010;
292 :  {high,med,low}<='h010;
293 :  {high,med,low}<='h010;
294 :  {high,med,low}<='h007;
295 :  {high,med,low}<='h007;
296 :  {high,med,low}<='h006;
297 :  {high,med,low}<='h006;
298 :  {high,med,low}<='h007;
299 :  {high,med,low}<='h007;
300 :  {high,med,low}<='h010;
301 :  {high,med,low}<='h010;
302 :  {high,med,low}<='h010;
303 :  {high,med,low}<='h010;
//20
304 :  {high,med,low}<='h000;
305 :  {high,med,low}<='h000;
306 :  {high,med,low}<='h007;
307 :  {high,med,low}<='h007;
308 :  {high,med,low}<='h006;
309 :  {high,med,low}<='h006;
310 :  {high,med,low}<='h007;
311 :  {high,med,low}<='h007;
312 :  {high,med,low}<='h010;
313 :  {high,med,low}<='h010;
314 :  {high,med,low}<='h020;
315 :  {high,med,low}<='h020;
316 :  {high,med,low}<='h030;
317 :  {high,med,low}<='h030;
318 :  {high,med,low}<='h040;
319 :  {high,med,low}<='h040;
//21
320 :  {high,med,low}<='h040;
321 :  {high,med,low}<='h040;
322 :  {high,med,low}<='h010;
323 :  {high,med,low}<='h010;
324 :  {high,med,low}<='h010;
325 :  {high,med,low}<='h010;
326 :  {high,med,low}<='h020;
327 :  {high,med,low}<='h030;
328 :  {high,med,low}<='h020;
329 :  {high,med,low}<='h020;
330 :  {high,med,low}<='h010;
331 :  {high,med,low}<='h000;
332 :  {high,med,low}<='h010;
333 :  {high,med,low}<='h010;
334 :  {high,med,low}<='h010;
335 :  {high,med,low}<='h010;
//22
336 :  {high,med,low}<='h000;
337 :  {high,med,low}<='h000;
338 :  {high,med,low}<='h000;
339 :  {high,med,low}<='h000;
340 :  {high,med,low}<='h000;
341 :  {high,med,low}<='h000;
342 :  {high,med,low}<='h000;
343 :  {high,med,low}<='h000;
344 :  {high,med,low}<='h000;
345 :  {high,med,low}<='h000;
346 :  {high,med,low}<='h000;
347 :  {high,med,low}<='h000;
348 :  {high,med,low}<='h030;
349 :  {high,med,low}<='h030;
350 :  {high,med,low}<='h050;
351 :  {high,med,low}<='h030;
//23
352 :  {high,med,low}<='h020;
353 :  {high,med,low}<='h020;
354 :  {high,med,low}<='h010;
355 :  {high,med,low}<='h010;
356 :  {high,med,low}<='h006;
357 :  {high,med,low}<='h010;
358 :  {high,med,low}<='h010;
359 :  {high,med,low}<='h020;
360 :  {high,med,low}<='h020;
361 :  {high,med,low}<='h020;
362 :  {high,med,low}<='h000;
363 :  {high,med,low}<='h000;
364 :  {high,med,low}<='h030;
365 :  {high,med,low}<='h030;
366 :  {high,med,low}<='h050;
367 :  {high,med,low}<='h030;
//24
368 :  {high,med,low}<='h020;
369 :  {high,med,low}<='h020;
370 :  {high,med,low}<='h010;
371 :  {high,med,low}<='h010;
372 :  {high,med,low}<='h005;
373 :  {high,med,low}<='h010;
374 :  {high,med,low}<='h010;
375 :  {high,med,low}<='h010;
376 :  {high,med,low}<='h010;
377 :  {high,med,low}<='h010;
378 :  {high,med,low}<='h000;
379 :  {high,med,low}<='h000;
380 :  {high,med,low}<='h030;
381 :  {high,med,low}<='h030;
382 :  {high,med,low}<='h050;
383 :  {high,med,low}<='h030;
//25
384 :  {high,med,low}<='h020;
385 :  {high,med,low}<='h020;
386 :  {high,med,low}<='h000;
387 :  {high,med,low}<='h000;
388 :  {high,med,low}<='h030;
389 :  {high,med,low}<='h050;
390 :  {high,med,low}<='h050;
391 :  {high,med,low}<='h050;
392 :  {high,med,low}<='h050;
393 :  {high,med,low}<='h060;
394 :  {high,med,low}<='h060;
395 :  {high,med,low}<='h060;
396 :  {high,med,low}<='h050;
397 :  {high,med,low}<='h040;
398 :  {high,med,low}<='h030;
399 :  {high,med,low}<='h030;
//26
400 :  {high,med,low}<='h030;
401 :  {high,med,low}<='h030;
402 :  {high,med,low}<='h030;
403 :  {high,med,low}<='h030;
404 :  {high,med,low}<='h030;
405 :  {high,med,low}<='h030;
406 :  {high,med,low}<='h030;
407 :  {high,med,low}<='h030;
408 :  {high,med,low}<='h000;
409 :  {high,med,low}<='h000;
410 :  {high,med,low}<='h000;
411 :  {high,med,low}<='h000;
412 :  {high,med,low}<='h030;
413 :  {high,med,low}<='h030;
414 :  {high,med,low}<='h050;
415 :  {high,med,low}<='h030;
//27
416 :  {high,med,low}<='h020;
417 :  {high,med,low}<='h020;
418 :  {high,med,low}<='h010;
419 :  {high,med,low}<='h010;
420 :  {high,med,low}<='h006;
421 :  {high,med,low}<='h010;
422 :  {high,med,low}<='h010;
423 :  {high,med,low}<='h002;
424 :  {high,med,low}<='h002;
425 :  {high,med,low}<='h002;
426 :  {high,med,low}<='h000;
427 :  {high,med,low}<='h000;
428 :  {high,med,low}<='h030;
429 :  {high,med,low}<='h030;
430 :  {high,med,low}<='h050;
431 :  {high,med,low}<='h030;
//28
432 :  {high,med,low}<='h020;
433 :  {high,med,low}<='h020;
434 :  {high,med,low}<='h010;
435 :  {high,med,low}<='h010;
436 :  {high,med,low}<='h006;
437 :  {high,med,low}<='h010;
438 :  {high,med,low}<='h010;
439 :  {high,med,low}<='h010;
440 :  {high,med,low}<='h010;
441 :  {high,med,low}<='h010;
442 :  {high,med,low}<='h000;
443 :  {high,med,low}<='h000;
444 :  {high,med,low}<='h010;
445 :  {high,med,low}<='h007;
446 :  {high,med,low}<='h006;
447 :  {high,med,low}<='h007;
//29
448 :  {high,med,low}<='h006;
449 :  {high,med,low}<='h006;
450 :  {high,med,low}<='h006;
451 :  {high,med,low}<='h006;
452 :  {high,med,low}<='h020;
453 :  {high,med,low}<='h020;
454 :  {high,med,low}<='h020;
455 :  {high,med,low}<='h020;
456 :  {high,med,low}<='h007;
457 :  {high,med,low}<='h007;
458 :  {high,med,low}<='h006;
459 :  {high,med,low}<='h006;
460 :  {high,med,low}<='h007;
461 :  {high,med,low}<='h000;
462 :  {high,med,low}<='h007;
463 :  {high,med,low}<='h007;
//30
464 :  {high,med,low}<='h007;
465 :  {high,med,low}<='h007;
466 :  {high,med,low}<='h010;
467 :  {high,med,low}<='h010;
468 :  {high,med,low}<='h010;
469 :  {high,med,low}<='h010;
470 :  {high,med,low}<='h010;
471 :  {high,med,low}<='h010;
472 :  {high,med,low}<='h010;
473 :  {high,med,low}<='h010;
474 :  {high,med,low}<='h010;
475 :  {high,med,low}<='h010;
476 :  {high,med,low}<='h000;
477 :  {high,med,low}<='h000;
478 :  {high,med,low}<='h000;
479 :  {high,med,low}<='h000;
//31
480 :  {high,med,low}<='h020;
481 :  {high,med,low}<='h020;
482 :  {high,med,low}<='h030;
483 :  {high,med,low}<='h030;
484 :  {high,med,low}<='h050;
485 :  {high,med,low}<='h050;
486 :  {high,med,low}<='h010;
487 :  {high,med,low}<='h010;
488 :  {high,med,low}<='h020;
489 :  {high,med,low}<='h020;
490 :  {high,med,low}<='h030;
491 :  {high,med,low}<='h030;
492 :  {high,med,low}<='h050;
493 :  {high,med,low}<='h050;
494 :  {high,med,low}<='h010;
495 :  {high,med,low}<='h010;
//32
496 :  {high,med,low}<='h020;
497 :  {high,med,low}<='h020;
498 :  {high,med,low}<='h030;
499 :  {high,med,low}<='h030;
500 :  {high,med,low}<='h050;
501 :  {high,med,low}<='h050;
502 :  {high,med,low}<='h060;
503 :  {high,med,low}<='h060;
504 :  {high,med,low}<='h020;
505 :  {high,med,low}<='h020;
506 :  {high,med,low}<='h030;
507 :  {high,med,low}<='h030;
508 :  {high,med,low}<='h006;
509 :  {high,med,low}<='h006;
510 :  {high,med,low}<='h010;
511 :  {high,med,low}<='h010;
//33
512 :  {high,med,low}<='h020;
513 :  {high,med,low}<='h020;
514 :  {high,med,low}<='h030;
515 :  {high,med,low}<='h030;
516 :  {high,med,low}<='h050;
517 :  {high,med,low}<='h050;
518 :  {high,med,low}<='h010;
519 :  {high,med,low}<='h010;
520 :  {high,med,low}<='h020;
521 :  {high,med,low}<='h020;
522 :  {high,med,low}<='h030;
523 :  {high,med,low}<='h030;
524 :  {high,med,low}<='h050;
525 :  {high,med,low}<='h050;
526 :  {high,med,low}<='h010;
527 :  {high,med,low}<='h010;
//34
528 :  {high,med,low}<='h020;
529 :  {high,med,low}<='h020;
530 :  {high,med,low}<='h030;
531 :  {high,med,low}<='h030;
532 :  {high,med,low}<='h050;
533 :  {high,med,low}<='h050;
534 :  {high,med,low}<='h060;
535 :  {high,med,low}<='h060;
536 :  {high,med,low}<='h020;
537 :  {high,med,low}<='h020;
538 :  {high,med,low}<='h030;
539 :  {high,med,low}<='h030;
540 :  {high,med,low}<='h000;
541 :  {high,med,low}<='h000;
542 :  {high,med,low}<='h010;
543 :  {high,med,low}<='h020;
//35
544 :  {high,med,low}<='h030;
545 :  {high,med,low}<='h030;
546 :  {high,med,low}<='h020;
547 :  {high,med,low}<='h010;
548 :  {high,med,low}<='h010;
549 :  {high,med,low}<='h010;
550 :  {high,med,low}<='h006;
551 :  {high,med,low}<='h007;
552 :  {high,med,low}<='h010;
553 :  {high,med,low}<='h010;
554 :  {high,med,low}<='h007;
555 :  {high,med,low}<='h006;
556 :  {high,med,low}<='h005;
557 :  {high,med,low}<='h005;
558 :  {high,med,low}<='h003;
559 :  {high,med,low}<='h005;
//36
560 :  {high,med,low}<='h006;
561 :  {high,med,low}<='h006;
562 :  {high,med,low}<='h007;
563 :  {high,med,low}<='h010;
564 :  {high,med,low}<='h007;
565 :  {high,med,low}<='h005;
566 :  {high,med,low}<='h005;
567 :  {high,med,low}<='h006;
568 :  {high,med,low}<='h005;
569 :  {high,med,low}<='h005;
570 :  {high,med,low}<='h005;
571 :  {high,med,low}<='h005;
572 :  {high,med,low}<='h003;
573 :  {high,med,low}<='h003;
574 :  {high,med,low}<='h005;
575 :  {high,med,low}<='h005;
//37
576 :  {high,med,low}<='h006;
577 :  {high,med,low}<='h006;
578 :  {high,med,low}<='h007;
579 :  {high,med,low}<='h010;
580 :  {high,med,low}<='h007;
581 :  {high,med,low}<='h007;
582 :  {high,med,low}<='h010;
583 :  {high,med,low}<='h020;
584 :  {high,med,low}<='h030;
585 :  {high,med,low}<='h030;
586 :  {high,med,low}<='h020;
587 :  {high,med,low}<='h010;
588 :  {high,med,low}<='h007;
589 :  {high,med,low}<='h007;
590 :  {high,med,low}<='h005;
591 :  {high,med,low}<='h000;
//38
592 :  {high,med,low}<='h005;
593 :  {high,med,low}<='h005;
594 :  {high,med,low}<='h005;
595 :  {high,med,low}<='h005;
596 :  {high,med,low}<='h000;
597 :  {high,med,low}<='h000;
598 :  {high,med,low}<='h000;
599 :  {high,med,low}<='h000;
600 :  {high,med,low}<='h000;
601 :  {high,med,low}<='h000;
602 :  {high,med,low}<='h000;
603 :  {high,med,low}<='h000;
604 :  {high,med,low}<='h000;
605 :  {high,med,low}<='h000;
606 :  {high,med,low}<='h010;
607 :  {high,med,low}<='h020;
//39
608 :  {high,med,low}<='h030;
609 :  {high,med,low}<='h030;
610 :  {high,med,low}<='h020;
611 :  {high,med,low}<='h010;
612 :  {high,med,low}<='h010;
613 :  {high,med,low}<='h010;
614 :  {high,med,low}<='h006;
615 :  {high,med,low}<='h007;
616 :  {high,med,low}<='h010;
617 :  {high,med,low}<='h010;
618 :  {high,med,low}<='h007;
619 :  {high,med,low}<='h006;
620 :  {high,med,low}<='h005;
621 :  {high,med,low}<='h005;
622 :  {high,med,low}<='h000;
623 :  {high,med,low}<='h005;
//40
624 :  {high,med,low}<='h006;
625 :  {high,med,low}<='h006;
626 :  {high,med,low}<='h007;
627 :  {high,med,low}<='h010;
628 :  {high,med,low}<='h007;
629 :  {high,med,low}<='h005;
630 :  {high,med,low}<='h005;
631 :  {high,med,low}<='h006;
632 :  {high,med,low}<='h005;
633 :  {high,med,low}<='h005;
634 :  {high,med,low}<='h000;
635 :  {high,med,low}<='h000;
636 :  {high,med,low}<='h006;
637 :  {high,med,low}<='h006;
638 :  {high,med,low}<='h006;
639 :  {high,med,low}<='h005;
//41
640 :  {high,med,low}<='h005;
641 :  {high,med,low}<='h005;
642 :  {high,med,low}<='h006;
643 :  {high,med,low}<='h006;
644 :  {high,med,low}<='h006;
645 :  {high,med,low}<='h010;
646 :  {high,med,low}<='h010;
647 :  {high,med,low}<='h010;
648 :  {high,med,low}<='h020;
649 :  {high,med,low}<='h020;
650 :  {high,med,low}<='h020;
651 :  {high,med,low}<='h030;
652 :  {high,med,low}<='h030;
653 :  {high,med,low}<='h030;
654 :  {high,med,low}<='h020;
655 :  {high,med,low}<='h020;
//42
656 :  {high,med,low}<='h010;
657 :  {high,med,low}<='h00;
658 :  {high,med,low}<='h010;
659 :  {high,med,low}<='h010;
660 :  {high,med,low}<='h010;
661 :  {high,med,low}<='h010;
662 :  {high,med,low}<='h010;
663 :  {high,med,low}<='h010;
664 :  {high,med,low}<='h000;
665 :  {high,med,low}<='h000;
666 :  {high,med,low}<='h000;
667 :  {high,med,low}<='h000;
668 :  {high,med,low}<='h000;
669 :  {high,med,low}<='h000;
670 :  {high,med,low}<='h000;
671 :  {high,med,low}<='h000;
//43
672 :  {high,med,low}<='h060;
673 :  {high,med,low}<='h060;
674 :  {high,med,low}<='h060;
675 :  {high,med,low}<='h060;
676 :  {high,med,low}<='h050;
677 :  {high,med,low}<='h050;
678 :  {high,med,low}<='h040;
679 :  {high,med,low}<='h040;
680 :  {high,med,low}<='h030;
681 :  {high,med,low}<='h030;
682 :  {high,med,low}<='h030;
683 :  {high,med,low}<='h030;
684 :  {high,med,low}<='h020;
685 :  {high,med,low}<='h030;
686 :  {high,med,low}<='h040;
687 :  {high,med,low}<='h040;
//44
688 :  {high,med,low}<='h040;
689 :  {high,med,low}<='h030;
690 :  {high,med,low}<='h020;
691 :  {high,med,low}<='h010;
692 :  {high,med,low}<='h010;
693 :  {high,med,low}<='h020;
694 :  {high,med,low}<='h030;
695 :  {high,med,low}<='h040;
696 :  {high,med,low}<='h040;
697 :  {high,med,low}<='h030;
698 :  {high,med,low}<='h020;
699 :  {high,med,low}<='h010;
700 :  {high,med,low}<='h010;
701 :  {high,med,low}<='h006;
702 :  {high,med,low}<='h007;
703 :  {high,med,low}<='h010;
//45
704 :  {high,med,low}<='h010;
705 :  {high,med,low}<='h007;
706 :  {high,med,low}<='h006;
707 :  {high,med,low}<='h005;
708 :  {high,med,low}<='h005;
709 :  {high,med,low}<='h005;
710 :  {high,med,low}<='h005;
711 :  {high,med,low}<='h005;
712 :  {high,med,low}<='h006;
713 :  {high,med,low}<='h006;
714 :  {high,med,low}<='h006;
715 :  {high,med,low}<='h010;
716 :  {high,med,low}<='h010;
717 :  {high,med,low}<='h010;
718 :  {high,med,low}<='h007;
719 :  {high,med,low}<='h007;
//46
720 :  {high,med,low}<='h007;
721 :  {high,med,low}<='h005;
722 :  {high,med,low}<='h005;
723 :  {high,med,low}<='h003;
724 :  {high,med,low}<='h003;
725 :  {high,med,low}<='h003;
726 :  {high,med,low}<='h003;
727 :  {high,med,low}<='h006;
728 :  {high,med,low}<='h006;
729 :  {high,med,low}<='h006;
730 :  {high,med,low}<='h006;
731 :  {high,med,low}<='h006;
732 :  {high,med,low}<='h006;
733 :  {high,med,low}<='h006;
734 :  {high,med,low}<='h006;
735 :  {high,med,low}<='h006;
//47
736 :  {high,med,low}<='h060;
737 :  {high,med,low}<='h060;
738 :  {high,med,low}<='h060;
739 :  {high,med,low}<='h060;
740 :  {high,med,low}<='h050;
741 :  {high,med,low}<='h050;
742 :  {high,med,low}<='h040;
743 :  {high,med,low}<='h040;
744 :  {high,med,low}<='h030;
745 :  {high,med,low}<='h030;
746 :  {high,med,low}<='h030;
747 :  {high,med,low}<='h030;
748 :  {high,med,low}<='h020;
749 :  {high,med,low}<='h030;
750 :  {high,med,low}<='h040;
751 :  {high,med,low}<='h040;
//48
752 :  {high,med,low}<='h040;
753 :  {high,med,low}<='h040;
754 :  {high,med,low}<='h040;
755 :  {high,med,low}<='h040;
756 :  {high,med,low}<='h030;
757 :  {high,med,low}<='h020;
758 :  {high,med,low}<='h030;
759 :  {high,med,low}<='h030;
760 :  {high,med,low}<='h030;
761 :  {high,med,low}<='h030;
762 :  {high,med,low}<='h030;
763 :  {high,med,low}<='h030;
764 :  {high,med,low}<='h000;
765 :  {high,med,low}<='h000;
766 :  {high,med,low}<='h000;
767 :  {high,med,low}<='h000;
//49
768 :  {high,med,low}<='h000;
769 :  {high,med,low}<='h000;
770 :  {high,med,low}<='h000;
771 :  {high,med,low}<='h000;
772 :  {high,med,low}<='h000;
773 :  {high,med,low}<='h000;
774 :  {high,med,low}<='h040;
775 :  {high,med,low}<='h040;
776 :  {high,med,low}<='h030;
777 :  {high,med,low}<='h030;
778 :  {high,med,low}<='h020;
779 :  {high,med,low}<='h020;
780 :  {high,med,low}<='h010;
781 :  {high,med,low}<='h010;
782 :  {high,med,low}<='h010;
783 :  {high,med,low}<='h010;
//50
784 :  {high,med,low}<='h000;
785 :  {high,med,low}<='h000;
786 :  {high,med,low}<='h000;
787 :  {high,med,low}<='h000;
788 :  {high,med,low}<='h000;
789 :  {high,med,low}<='h000;
790 :  {high,med,low}<='h000;
791 :  {high,med,low}<='h000;
792 :  {high,med,low}<='h000;
793 :  {high,med,low}<='h000;
794 :  {high,med,low}<='h000;
795 :  {high,med,low}<='h000;
796 :  {high,med,low}<='h030;
797 :  {high,med,low}<='h030;
798 :  {high,med,low}<='h050;
799 :  {high,med,low}<='h030;
//51
800 :  {high,med,low}<='h020;
801 :  {high,med,low}<='h020;
802 :  {high,med,low}<='h010;
803 :  {high,med,low}<='h010;
804 :  {high,med,low}<='h006;
805 :  {high,med,low}<='h010;
806 :  {high,med,low}<='h010;
807 :  {high,med,low}<='h020;
808 :  {high,med,low}<='h020;
809 :  {high,med,low}<='h020;
810 :  {high,med,low}<='h000;
811 :  {high,med,low}<='h000;
812 :  {high,med,low}<='h030;
813 :  {high,med,low}<='h030;
814 :  {high,med,low}<='h050;
815 :  {high,med,low}<='h030;
//52
816 :  {high,med,low}<='h020;
817 :  {high,med,low}<='h020;
818 :  {high,med,low}<='h010;
819 :  {high,med,low}<='h010;
820 :  {high,med,low}<='h006;
821 :  {high,med,low}<='h010;
822 :  {high,med,low}<='h010;
823 :  {high,med,low}<='h010;
824 :  {high,med,low}<='h010;
825 :  {high,med,low}<='h010;
826 :  {high,med,low}<='h000;
827 :  {high,med,low}<='h000;
828 :  {high,med,low}<='h030;
829 :  {high,med,low}<='h030;
830 :  {high,med,low}<='h050;
831 :  {high,med,low}<='h030;
//53
832 :  {high,med,low}<='h020;
833 :  {high,med,low}<='h020;
834 :  {high,med,low}<='h000;
835 :  {high,med,low}<='h000;
836 :  {high,med,low}<='h030;
837 :  {high,med,low}<='h050;
838 :  {high,med,low}<='h050;
839 :  {high,med,low}<='h050;
840 :  {high,med,low}<='h050;
841 :  {high,med,low}<='h060;
842 :  {high,med,low}<='h060;
843 :  {high,med,low}<='h060;
844 :  {high,med,low}<='h050;
845 :  {high,med,low}<='h040;
846 :  {high,med,low}<='h030;
847 :  {high,med,low}<='h030;
//54
848 :  {high,med,low}<='h030;
849 :  {high,med,low}<='h030;
850 :  {high,med,low}<='h030;
851 :  {high,med,low}<='h030;
852 :  {high,med,low}<='h030;
853 :  {high,med,low}<='h030;
854 :  {high,med,low}<='h030;
855 :  {high,med,low}<='h030;
856 :  {high,med,low}<='h000;
857 :  {high,med,low}<='h000;
858 :  {high,med,low}<='h000;
859 :  {high,med,low}<='h000;
860 :  {high,med,low}<='h030;
861 :  {high,med,low}<='h030;
862 :  {high,med,low}<='h050;
863 :  {high,med,low}<='h030;
//55
864 :  {high,med,low}<='h020;
865 :  {high,med,low}<='h020;
866 :  {high,med,low}<='h010;
867 :  {high,med,low}<='h010;
868 :  {high,med,low}<='h006;
869 :  {high,med,low}<='h010;
870 :  {high,med,low}<='h010;
871 :  {high,med,low}<='h020;
872 :  {high,med,low}<='h020;
873 :  {high,med,low}<='h020;
874 :  {high,med,low}<='h000;
875 :  {high,med,low}<='h000;
876 :  {high,med,low}<='h030;
877 :  {high,med,low}<='h030;
878 :  {high,med,low}<='h050;
879 :  {high,med,low}<='h030;
//56
880 :  {high,med,low}<='h020;
881 :  {high,med,low}<='h020;
882 :  {high,med,low}<='h010;
883 :  {high,med,low}<='h010;
884 :  {high,med,low}<='h006;
885 :  {high,med,low}<='h010;
886 :  {high,med,low}<='h010;
887 :  {high,med,low}<='h010;
888 :  {high,med,low}<='h010;
889 :  {high,med,low}<='h010;
890 :  {high,med,low}<='h000;
891 :  {high,med,low}<='h000;
892 :  {high,med,low}<='h010;
893 :  {high,med,low}<='h070;
894 :  {high,med,low}<='h060;
895 :  {high,med,low}<='h070;
//57
896 :  {high,med,low}<='h006;
897 :  {high,med,low}<='h006;
898 :  {high,med,low}<='h006;
899 :  {high,med,low}<='h006;
900 :  {high,med,low}<='h020;
901 :  {high,med,low}<='h020;
902 :  {high,med,low}<='h020;
903 :  {high,med,low}<='h020;
904 :  {high,med,low}<='h007;
905 :  {high,med,low}<='h007;
906 :  {high,med,low}<='h005;
907 :  {high,med,low}<='h005;
908 :  {high,med,low}<='h003;
909 :  {high,med,low}<='h003;
910 :  {high,med,low}<='h007;
911 :  {high,med,low}<='h007;
//58
912 :  {high,med,low}<='h007;
913 :  {high,med,low}<='h007;
914 :  {high,med,low}<='h010;
915 :  {high,med,low}<='h010;
916 :  {high,med,low}<='h010;
917 :  {high,med,low}<='h010;
918 :  {high,med,low}<='h010;
919 :  {high,med,low}<='h010;
920 :  {high,med,low}<='h000;
921 :  {high,med,low}<='h000;
922 :  {high,med,low}<='h000;
923 :  {high,med,low}<='h000;
924 :  {high,med,low}<='h000;
925 :  {high,med,low}<='h000;
926 :  {high,med,low}<='h000;
927 :  {high,med,low}<='h000;
//59
928 :  {high,med,low}<='h000;
929 :  {high,med,low}<='h000;
930 :  {high,med,low}<='h050;
931 :  {high,med,low}<='h050;
932 :  {high,med,low}<='h030;
933 :  {high,med,low}<='h020;
934 :  {high,med,low}<='h010;
935 :  {high,med,low}<='h020;
936 :  {high,med,low}<='h000;
937 :  {high,med,low}<='h020;
938 :  {high,med,low}<='h020;
939 :  {high,med,low}<='h020;
940 :  {high,med,low}<='h020;
941 :  {high,med,low}<='h020;
942 :  {high,med,low}<='h020;
943 :  {high,med,low}<='h020;
//60
944 :  {high,med,low}<='h000;
945 :  {high,med,low}<='h000;
946 :  {high,med,low}<='h050;
947 :  {high,med,low}<='h050;
948 :  {high,med,low}<='h030;
949 :  {high,med,low}<='h020;
950 :  {high,med,low}<='h010;
951 :  {high,med,low}<='h020;
952 :  {high,med,low}<='h000;
953 :  {high,med,low}<='h020;
954 :  {high,med,low}<='h020;
955 :  {high,med,low}<='h020;
956 :  {high,med,low}<='h020;
957 :  {high,med,low}<='h020;
958 :  {high,med,low}<='h020;
959 :  {high,med,low}<='h020;
//61
960 :  {high,med,low}<='h000;
961 :  {high,med,low}<='h000;
962 :  {high,med,low}<='h050;
963 :  {high,med,low}<='h050;
964 :  {high,med,low}<='h030;
965 :  {high,med,low}<='h020;
966 :  {high,med,low}<='h010;
967 :  {high,med,low}<='h020;
968 :  {high,med,low}<='h020;
969 :  {high,med,low}<='h020;
970 :  {high,med,low}<='h020;
971 :  {high,med,low}<='h020;
972 :  {high,med,low}<='h020;
973 :  {high,med,low}<='h020;
974 :  {high,med,low}<='h020;
975 :  {high,med,low}<='h020;
//62
976 :  {high,med,low}<='h000;
977 :  {high,med,low}<='h000;
978 :  {high,med,low}<='h060;
979 :  {high,med,low}<='h060;
980 :  {high,med,low}<='h050;
981 :  {high,med,low}<='h040;
982 :  {high,med,low}<='h040;
983 :  {high,med,low}<='h050;
984 :  {high,med,low}<='h050;
985 :  {high,med,low}<='h050;
986 :  {high,med,low}<='h050;
987 :  {high,med,low}<='h050;
988 :  {high,med,low}<='h050;
989 :  {high,med,low}<='h050;
990 :  {high,med,low}<='h050;
991 :  {high,med,low}<='h050;
//63
992 :  {high,med,low}<='h000;
993 :  {high,med,low}<='h000;
994 :  {high,med,low}<='h050;
995 :  {high,med,low}<='h050;
996 :  {high,med,low}<='h030;
997 :  {high,med,low}<='h020;
998 :  {high,med,low}<='h010;
999 :  {high,med,low}<='h020;
1000 :  {high,med,low}<='h000;
1001 :  {high,med,low}<='h020;
1002 :  {high,med,low}<='h020;
1003 :  {high,med,low}<='h020;
1004 :  {high,med,low}<='h020;
1005 :  {high,med,low}<='h020;
1006 :  {high,med,low}<='h020;
1007 :  {high,med,low}<='h020;
//64
1008 :  {high,med,low}<='h000;
1009 :  {high,med,low}<='h000;
1010 :  {high,med,low}<='h050;
1011 :  {high,med,low}<='h050;
1012 :  {high,med,low}<='h030;
1013 :  {high,med,low}<='h020;
1014 :  {high,med,low}<='h010;
1015 :  {high,med,low}<='h020;
1016 :  {high,med,low}<='h000;
1017 :  {high,med,low}<='h020;
1018 :  {high,med,low}<='h020;
1019 :  {high,med,low}<='h020;
1020 :  {high,med,low}<='h020;
1021 :  {high,med,low}<='h020;
1022 :  {high,med,low}<='h020;
1023 :  {high,med,low}<='h020;
//65
1024 :  {high,med,low}<='h000;
1025 :  {high,med,low}<='h000;
1026 :  {high,med,low}<='h050;
1027 :  {high,med,low}<='h050;
1028 :  {high,med,low}<='h030;
1029 :  {high,med,low}<='h020;
1030 :  {high,med,low}<='h010;
1031 :  {high,med,low}<='h020;
1032 :  {high,med,low}<='h020;
1033 :  {high,med,low}<='h020;
1034 :  {high,med,low}<='h010;
1035 :  {high,med,low}<='h020;
1036 :  {high,med,low}<='h030;
1037 :  {high,med,low}<='h030;
1038 :  {high,med,low}<='h040;
1039 :  {high,med,low}<='h040;
//66
1040 :  {high,med,low}<='h020;
1041 :  {high,med,low}<='h000;
1042 :  {high,med,low}<='h020;
1043 :  {high,med,low}<='h020;
1044 :  {high,med,low}<='h020;
1045 :  {high,med,low}<='h020;
1046 :  {high,med,low}<='h020;
1047 :  {high,med,low}<='h020;
1048 :  {high,med,low}<='h000;
1049 :  {high,med,low}<='h000;
1050 :  {high,med,low}<='h000;
1051 :  {high,med,low}<='h000;
1052 :  {high,med,low}<='h000;
1053 :  {high,med,low}<='h000;
1054 :  {high,med,low}<='h000;
1055 :  {high,med,low}<='h000;
//67
1056 :  {high,med,low}<='h200;
1057 :  {high,med,low}<='h200;
1058 :  {high,med,low}<='h300;
1059 :  {high,med,low}<='h300;
1060 :  {high,med,low}<='h500;
1061 :  {high,med,low}<='h500;
1062 :  {high,med,low}<='h100;
1063 :  {high,med,low}<='h100;
1064 :  {high,med,low}<='h200;
1065 :  {high,med,low}<='h200;
1066 :  {high,med,low}<='h300;
1067 :  {high,med,low}<='h300;
1068 :  {high,med,low}<='h500;
1069 :  {high,med,low}<='h500;
1070 :  {high,med,low}<='h100;
1071 :  {high,med,low}<='h100;
//68
1072 :  {high,med,low}<='h200;
1073 :  {high,med,low}<='h200;
1074 :  {high,med,low}<='h300;
1075 :  {high,med,low}<='h300;
1076 :  {high,med,low}<='h500;
1077 :  {high,med,low}<='h500;
1078 :  {high,med,low}<='h100;
1079 :  {high,med,low}<='h100;
1080 :  {high,med,low}<='h200;
1081 :  {high,med,low}<='h200;
1082 :  {high,med,low}<='h300;
1083 :  {high,med,low}<='h300;
1084 :  {high,med,low}<='h500;
1085 :  {high,med,low}<='h500;
1086 :  {high,med,low}<='h100;
1087 :  {high,med,low}<='h100;
//69
1088 :  {high,med,low}<='h200;
1089 :  {high,med,low}<='h200;
1090 :  {high,med,low}<='h300;
1091 :  {high,med,low}<='h300;
1092 :  {high,med,low}<='h500;
1093 :  {high,med,low}<='h500;
1094 :  {high,med,low}<='h100;
1095 :  {high,med,low}<='h100;
1096 :  {high,med,low}<='h200;
1097 :  {high,med,low}<='h200;
1098 :  {high,med,low}<='h300;
1099 :  {high,med,low}<='h300;
1100 :  {high,med,low}<='h500;
1101 :  {high,med,low}<='h500;
1102 :  {high,med,low}<='h100;
1103 :  {high,med,low}<='h100;
//70
1104 :  {high,med,low}<='h200;
1105 :  {high,med,low}<='h200;
1106 :  {high,med,low}<='h300;
1107 :  {high,med,low}<='h300;
1108 :  {high,med,low}<='h500;
1109 :  {high,med,low}<='h500;
1110 :  {high,med,low}<='h100;
1111 :  {high,med,low}<='h100;
1112 :  {high,med,low}<='h200;
1113 :  {high,med,low}<='h200;
1114 :  {high,med,low}<='h300;
1115 :  {high,med,low}<='h300;
1116 :  {high,med,low}<='h003;
1117 :  {high,med,low}<='h003;
1118 :  {high,med,low}<='h005;
1119 :  {high,med,low}<='h005;
//71
1120 :  {high,med,low}<='h006;
1121 :  {high,med,low}<='h006;
1122 :  {high,med,low}<='h006;
1123 :  {high,med,low}<='h006;
1124 :  {high,med,low}<='h010;
1125 :  {high,med,low}<='h010;
1126 :  {high,med,low}<='h020;
1127 :  {high,med,low}<='h020;
1128 :  {high,med,low}<='h020;
1129 :  {high,med,low}<='h020;
1130 :  {high,med,low}<='h010;
1131 :  {high,med,low}<='h010;
1132 :  {high,med,low}<='h005;
1133 :  {high,med,low}<='h005;
1134 :  {high,med,low}<='h004;
1135 :  {high,med,low}<='h004;
//72
1136 :  {high,med,low}<='h003;
1137 :  {high,med,low}<='h003;
1138 :  {high,med,low}<='h005;
1139 :  {high,med,low}<='h005;
1140 :  {high,med,low}<='h010;
1141 :  {high,med,low}<='h010;
1142 :  {high,med,low}<='h010;
1143 :  {high,med,low}<='h010;
1144 :  {high,med,low}<='h000;
1145 :  {high,med,low}<='h000;
1146 :  {high,med,low}<='h000;
1147 :  {high,med,low}<='h000;
1148 :  {high,med,low}<='h010;
1149 :  {high,med,low}<='h010;
1150 :  {high,med,low}<='h007;
1151 :  {high,med,low}<='h007;
//73
1152 :  {high,med,low}<='h006;
1153 :  {high,med,low}<='h006;
1154 :  {high,med,low}<='h006;
1155 :  {high,med,low}<='h006;
1156 :  {high,med,low}<='h010;
1157 :  {high,med,low}<='h010;
1158 :  {high,med,low}<='h010;
1159 :  {high,med,low}<='h010;
1160 :  {high,med,low}<='h007;
1161 :  {high,med,low}<='h007;
1162 :  {high,med,low}<='h005;
1163 :  {high,med,low}<='h005;
1164 :  {high,med,low}<='h005;
1165 :  {high,med,low}<='h000;
1166 :  {high,med,low}<='h005;
1167 :  {high,med,low}<='h005;
//74
1168 :  {high,med,low}<='h005;
1169 :  {high,med,low}<='h005;
1170 :  {high,med,low}<='h005;
1171 :  {high,med,low}<='h005;
1172 :  {high,med,low}<='h000;
1173 :  {high,med,low}<='h000;
1174 :  {high,med,low}<='h000;
1175 :  {high,med,low}<='h000;
1176 :  {high,med,low}<='h000;
1177 :  {high,med,low}<='h000;
1178 :  {high,med,low}<='h000;
1179 :  {high,med,low}<='h000;
1180 :  {high,med,low}<='h003;
1181 :  {high,med,low}<='h003;
1182 :  {high,med,low}<='h005;
1183 :  {high,med,low}<='h005;
//75
1184 :  {high,med,low}<='h006;
1185 :  {high,med,low}<='h006;
1186 :  {high,med,low}<='h006;
1187 :  {high,med,low}<='h006;
1188 :  {high,med,low}<='h010;
1189 :  {high,med,low}<='h010;
1190 :  {high,med,low}<='h020;
1191 :  {high,med,low}<='h020;
1192 :  {high,med,low}<='h020;
1193 :  {high,med,low}<='h020;
1194 :  {high,med,low}<='h010;
1195 :  {high,med,low}<='h010;
1196 :  {high,med,low}<='h005;
1197 :  {high,med,low}<='h005;
1198 :  {high,med,low}<='h004;
1199 :  {high,med,low}<='h004;
//76
1200 :  {high,med,low}<='h003;
1201 :  {high,med,low}<='h003;
1202 :  {high,med,low}<='h005;
1203 :  {high,med,low}<='h005;
1204 :  {high,med,low}<='h007;
1205 :  {high,med,low}<='h007;
1206 :  {high,med,low}<='h010;
1207 :  {high,med,low}<='h010;
1208 :  {high,med,low}<='h000;
1209 :  {high,med,low}<='h000;
1210 :  {high,med,low}<='h000;
1211 :  {high,med,low}<='h000;
1212 :  {high,med,low}<='h010;
1213 :  {high,med,low}<='h010;
1214 :  {high,med,low}<='h007;
1215 :  {high,med,low}<='h007;
//77
1216 :  {high,med,low}<='h006;
1217 :  {high,med,low}<='h006;
1218 :  {high,med,low}<='h006;
1219 :  {high,med,low}<='h006;
1220 :  {high,med,low}<='h010;
1221 :  {high,med,low}<='h010;
1222 :  {high,med,low}<='h010;
1223 :  {high,med,low}<='h010;
1224 :  {high,med,low}<='h007;
1225 :  {high,med,low}<='h007;
1226 :  {high,med,low}<='h005;
1227 :  {high,med,low}<='h005;
1228 :  {high,med,low}<='h005;
1229 :  {high,med,low}<='h005;
1230 :  {high,med,low}<='h006;
1231 :  {high,med,low}<='h006;
//78
1232 :  {high,med,low}<='h006;
1233 :  {high,med,low}<='h006;
1234 :  {high,med,low}<='h006;
1235 :  {high,med,low}<='h006;
1236 :  {high,med,low}<='h000;
1237 :  {high,med,low}<='h000;
1238 :  {high,med,low}<='h000;
1239 :  {high,med,low}<='h000;
1240 :  {high,med,low}<='h000;
1241 :  {high,med,low}<='h000;
1242 :  {high,med,low}<='h000;
1243 :  {high,med,low}<='h000;
1244 :  {high,med,low}<='h030;
1245 :  {high,med,low}<='h030;
1246 :  {high,med,low}<='h050;
1247 :  {high,med,low}<='h030;
//79
1248 :  {high,med,low}<='h020;
1249 :  {high,med,low}<='h020;
1250 :  {high,med,low}<='h010;
1251 :  {high,med,low}<='h010;
1252 :  {high,med,low}<='h006;
1253 :  {high,med,low}<='h010;
1254 :  {high,med,low}<='h010;
1255 :  {high,med,low}<='h020;
1256 :  {high,med,low}<='h020;
1257 :  {high,med,low}<='h020;
1258 :  {high,med,low}<='h000;
1259 :  {high,med,low}<='h000;
1260 :  {high,med,low}<='h030;
1261 :  {high,med,low}<='h030;
1262 :  {high,med,low}<='h050;
1263 :  {high,med,low}<='h030;
//80
1264 :  {high,med,low}<='h020;
1265 :  {high,med,low}<='h020;
1266 :  {high,med,low}<='h010;
1267 :  {high,med,low}<='h010;
1268 :  {high,med,low}<='h005;
1269 :  {high,med,low}<='h010;
1270 :  {high,med,low}<='h000;
1271 :  {high,med,low}<='h010;
1272 :  {high,med,low}<='h010;
1273 :  {high,med,low}<='h010;
1274 :  {high,med,low}<='h000;
1275 :  {high,med,low}<='h000;
1276 :  {high,med,low}<='h030;
1277 :  {high,med,low}<='h030;
1278 :  {high,med,low}<='h050;
1279 :  {high,med,low}<='h030;
//81
1280 :  {high,med,low}<='h020;
1281 :  {high,med,low}<='h020;
1282 :  {high,med,low}<='h000;
1283 :  {high,med,low}<='h000;
1284 :  {high,med,low}<='h030;
1285 :  {high,med,low}<='h050;
1286 :  {high,med,low}<='h050;
1287 :  {high,med,low}<='h050;
1288 :  {high,med,low}<='h050;
1289 :  {high,med,low}<='h060;
1290 :  {high,med,low}<='h060;
1291 :  {high,med,low}<='h060;
1292 :  {high,med,low}<='h050;
1293 :  {high,med,low}<='h040;
1294 :  {high,med,low}<='h030;
1295 :  {high,med,low}<='h030;
//82
1296 :  {high,med,low}<='h030;
1297 :  {high,med,low}<='h030;
1298 :  {high,med,low}<='h030;
1299 :  {high,med,low}<='h030;
1300 :  {high,med,low}<='h030;
1301 :  {high,med,low}<='h030;
1302 :  {high,med,low}<='h030;
1303 :  {high,med,low}<='h030;
1304 :  {high,med,low}<='h000;
1305 :  {high,med,low}<='h000;
1306 :  {high,med,low}<='h000;
1307 :  {high,med,low}<='h000;
1308 :  {high,med,low}<='h030;
1309 :  {high,med,low}<='h030;
1310 :  {high,med,low}<='h050;
1311 :  {high,med,low}<='h030;
//83
1312 :  {high,med,low}<='h020;
1313 :  {high,med,low}<='h020;
1314 :  {high,med,low}<='h010;
1315 :  {high,med,low}<='h010;
1316 :  {high,med,low}<='h006;
1317 :  {high,med,low}<='h010;
1318 :  {high,med,low}<='h010;
1319 :  {high,med,low}<='h020;
1320 :  {high,med,low}<='h020;
1321 :  {high,med,low}<='h020;
1322 :  {high,med,low}<='h000;
1323 :  {high,med,low}<='h000;
1324 :  {high,med,low}<='h030;
1325 :  {high,med,low}<='h030;
1326 :  {high,med,low}<='h050;
1327 :  {high,med,low}<='h030;
//84
1328 :  {high,med,low}<='h020;
1329 :  {high,med,low}<='h020;
1330 :  {high,med,low}<='h010;
1331 :  {high,med,low}<='h010;
1332 :  {high,med,low}<='h006;
1333 :  {high,med,low}<='h010;
1334 :  {high,med,low}<='h000;
1335 :  {high,med,low}<='h010;
1336 :  {high,med,low}<='h010;
1337 :  {high,med,low}<='h010;
1338 :  {high,med,low}<='h000;
1339 :  {high,med,low}<='h000;
1340 :  {high,med,low}<='h010;
1341 :  {high,med,low}<='h007;
1342 :  {high,med,low}<='h006;
1343 :  {high,med,low}<='h007;
//85
1344 :  {high,med,low}<='h006;
1345 :  {high,med,low}<='h006;
1346 :  {high,med,low}<='h000;
1347 :  {high,med,low}<='h006;
1348 :  {high,med,low}<='h020;
1349 :  {high,med,low}<='h020;
1350 :  {high,med,low}<='h020;
1351 :  {high,med,low}<='h020;
1352 :  {high,med,low}<='h007;
1353 :  {high,med,low}<='h007;
1354 :  {high,med,low}<='h006;
1355 :  {high,med,low}<='h006;
1356 :  {high,med,low}<='h007;
1357 :  {high,med,low}<='h007;
1358 :  {high,med,low}<='h007;
1359 :  {high,med,low}<='h000;
//86
1360 :  {high,med,low}<='h007;
1361 :  {high,med,low}<='h007;
1362 :  {high,med,low}<='h010;
1363 :  {high,med,low}<='h010;
1364 :  {high,med,low}<='h010;
1365 :  {high,med,low}<='h010;
1366 :  {high,med,low}<='h010;
1367 :  {high,med,low}<='h010;
1368 :  {high,med,low}<='h000;
1369 :  {high,med,low}<='h000;
1370 :  {high,med,low}<='h000;
1371 :  {high,med,low}<='h000;
1372 :  {high,med,low}<='h000;
1373 :  {high,med,low}<='h000;
1374 :  {high,med,low}<='h000;
1375 :  {high,med,low}<='h000;
//87
1376 :  {high,med,low}<='h006;
1377 :  {high,med,low}<='h006;
1378 :  {high,med,low}<='h006;
1379 :  {high,med,low}<='h000;
1380 :  {high,med,low}<='h006;
1381 :  {high,med,low}<='h007;
1382 :  {high,med,low}<='h010;
1383 :  {high,med,low}<='h010;
1384 :  {high,med,low}<='h020;
1385 :  {high,med,low}<='h020;
1386 :  {high,med,low}<='h020;
1387 :  {high,med,low}<='h020;
1388 :  {high,med,low}<='h030;
1389 :  {high,med,low}<='h030;
1390 :  {high,med,low}<='h010;
1391 :  {high,med,low}<='h000;
//88
1392 :  {high,med,low}<='h010;
1393 :  {high,med,low}<='h010;
1394 :  {high,med,low}<='h010;
1395 :  {high,med,low}<='h010;
1396 :  {high,med,low}<='h030;
1397 :  {high,med,low}<='h020;
1398 :  {high,med,low}<='h010;
1399 :  {high,med,low}<='h010;
1400 :  {high,med,low}<='h020;
1401 :  {high,med,low}<='h020;
1402 :  {high,med,low}<='h020;
1403 :  {high,med,low}<='h020;
1404 :  {high,med,low}<='h050;
1405 :  {high,med,low}<='h050;
1406 :  {high,med,low}<='h030;
1407 :  {high,med,low}<='h030;
//89
1408 :  {high,med,low}<='h030;
1409 :  {high,med,low}<='h030;
1410 :  {high,med,low}<='h030;
1411 :  {high,med,low}<='h030;
1412 :  {high,med,low}<='h010;
1413 :  {high,med,low}<='h010;
1414 :  {high,med,low}<='h005;
1415 :  {high,med,low}<='h005;
1416 :  {high,med,low}<='h006;
1417 :  {high,med,low}<='h006;
1418 :  {high,med,low}<='h006;
1419 :  {high,med,low}<='h006;
1420 :  {high,med,low}<='h005;
1421 :  {high,med,low}<='h005;
1422 :  {high,med,low}<='h004;
1423 :  {high,med,low}<='h004;
//90
1424 :  {high,med,low}<='h005;
1425 :  {high,med,low}<='h005;
1426 :  {high,med,low}<='h005;
1427 :  {high,med,low}<='h005;
1428 :  {high,med,low}<='h005;
1429 :  {high,med,low}<='h005;
1430 :  {high,med,low}<='h005;
1431 :  {high,med,low}<='h005;
1432 :  {high,med,low}<='h000;
1433 :  {high,med,low}<='h000;
1434 :  {high,med,low}<='h000;
1435 :  {high,med,low}<='h000;
1436 :  {high,med,low}<='h000;
1437 :  {high,med,low}<='h000;
1438 :  {high,med,low}<='h000;
1439 :  {high,med,low}<='h000;
//91
1440 :  {high,med,low}<='h006;
1441 :  {high,med,low}<='h006;
1442 :  {high,med,low}<='h006;
1443 :  {high,med,low}<='h000;
1444 :  {high,med,low}<='h006;
1445 :  {high,med,low}<='h007;
1446 :  {high,med,low}<='h010;
1447 :  {high,med,low}<='h010;
1448 :  {high,med,low}<='h020;
1449 :  {high,med,low}<='h020;
1450 :  {high,med,low}<='h020;
1451 :  {high,med,low}<='h020;
1452 :  {high,med,low}<='h030;
1453 :  {high,med,low}<='h030;
1454 :  {high,med,low}<='h010;
1455 :  {high,med,low}<='h010;
//92
1456 :  {high,med,low}<='h010;
1457 :  {high,med,low}<='h010;
1458 :  {high,med,low}<='h010;
1459 :  {high,med,low}<='h010;
1460 :  {high,med,low}<='h030;
1461 :  {high,med,low}<='h020;
1462 :  {high,med,low}<='h010;
1463 :  {high,med,low}<='h010;
1464 :  {high,med,low}<='h020;
1465 :  {high,med,low}<='h020;
1466 :  {high,med,low}<='h020;
1467 :  {high,med,low}<='h020;
1468 :  {high,med,low}<='h050;
1469 :  {high,med,low}<='h050;
1470 :  {high,med,low}<='h030;
1471 :  {high,med,low}<='h030;
//93
1472 :  {high,med,low}<='h060;
1473 :  {high,med,low}<='h060;
1474 :  {high,med,low}<='h060;
1475 :  {high,med,low}<='h060;
1476 :  {high,med,low}<='h060;
1477 :  {high,med,low}<='h060;
1478 :  {high,med,low}<='h030;
1479 :  {high,med,low}<='h030;
1480 :  {high,med,low}<='h020;
1481 :  {high,med,low}<='h020;
1482 :  {high,med,low}<='h020;
1483 :  {high,med,low}<='h020;
1484 :  {high,med,low}<='h020;
1485 :  {high,med,low}<='h020;
1486 :  {high,med,low}<='h010;
1487 :  {high,med,low}<='h020;
//94
1488 :  {high,med,low}<='h030;
1489 :  {high,med,low}<='h030;
1490 :  {high,med,low}<='h030;
1491 :  {high,med,low}<='h030;
1492 :  {high,med,low}<='h030;
1493 :  {high,med,low}<='h030;
1494 :  {high,med,low}<='h020;
1495 :  {high,med,low}<='h010;
1496 :  {high,med,low}<='h010;
1497 :  {high,med,low}<='h010;
1498 :  {high,med,low}<='h010;
1499 :  {high,med,low}<='h010;
1500 :  {high,med,low}<='h010;
1501 :  {high,med,low}<='h010;
1502 :  {high,med,low}<='h010;
1503 :  {high,med,low}<='h010;
//baba is you bgm
//0: {high,med,low}<='h005;
//1: {high,med,low}<='h000;
//2: {high,med,low}<='h000;
//3: {high,med,low}<='h000;
//4: {high,med,low}<='h000;
//5: {high,med,low}<='h000;
//6: {high,med,low}<='h000;
//7: {high,med,low}<='h000;
//8: {high,med,low}<='h000;
//9: {high,med,low}<='h000;
//10: {high,med,low}<='h000;
//11: {high,med,low}<='h000;
//12: {high,med,low}<='h000;
//13: {high,med,low}<='h000;
//14: {high,med,low}<='h004;
//15: {high,med,low}<='h000;
//16: {high,med,low}<='h000;
//17: {high,med,low}<='h000;
//18: {high,med,low}<='h000;
//19: {high,med,low}<='h000;
//20: {high,med,low}<='h000;
//21: {high,med,low}<='h000;
//22: {high,med,low}<='h000;
//23: {high,med,low}<='h000;
//24: {high,med,low}<='h000;
//25: {high,med,low}<='h000;
//26: {high,med,low}<='h000;
//27: {high,med,low}<='h000;
//28: {high,med,low}<='h002;
//29: {high,med,low}<='h002;
//30: {high,med,low}<='h000;

default: {high,med,low}<='h000;
    endcase
end
//led7s u1(high,high_7s);
//led7s u2(med,med_7s);
//led7s u3(low,low_7s);
endmodule